module sub(input [15:0] a, b, input cin, output [15:0] s, output cout);
	
	
	add a1 (a, ~b, cin, s, cout);
	
	


endmodule

